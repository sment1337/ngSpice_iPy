* This circuit contains only Berkeley SPICE3 components.
*
* The circuit is an AC coupled transistor amplifier with
* a sinewave input at node "1", a gain of approximately -3.9, * and output on node "coll".
*
.tran 1e-5 2e-3
*.dc vcc 0 15 0.1
*
vcc vcc 0 12.0
vin 1 0 0.0 ac 1.0 sin(0 1 1k)
ccouple 1 base 2.8300000000000002e-08
rbias1 vcc base 100k
rbias2 base 0 20000.0
q1 coll base emit generic
rcollector vcc coll 3.9k
remitter emit 0 200.0
*
.model generic npn
*.print dc coll
.print tran coll
* 
.end
